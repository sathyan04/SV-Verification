module half_adder(variables ha);
  assign {ha.carry,ha.sum}=a+b;
endmodule
