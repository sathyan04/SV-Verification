module half_adder(variables ha);
  assign {ha.cout,ha.sum}=a+b;
endmodule
